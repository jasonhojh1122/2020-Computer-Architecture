/*
ALU ALU(
    .data1_i    (),
    .data2_i    (),
    .ALUCtrl_i  (),
    .data_o     (),
    .Zero_o     ()
);
*/

module ALU
(
    data1_i,
    data2_i,
    ALUCtrl_i,
    data_o,
    Zero
);




endmodule